----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date: 07/23/2025 01:56:58 PM
-- Design Name: 
-- Module Name: data_memory - Behavioral
-- Project Name: 
-- Target Devices: 
-- Tool Versions: 
-- Description: 
-- 
-- Dependencies: 
-- 
-- Revision:
-- Revision 0.01 - File Created
-- Additional Comments:
-- 
----------------------------------------------------------------------------------


library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx leaf cells in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity data_memory is
    Port ( clk : in STD_LOGIC;
           wr_en : in STD_LOGIC;
           addr : in STD_LOGIC_VECTOR (7 downto 0);
           wr_data : in STD_LOGIC_VECTOR (31 downto 0);
           rd_data : out STD_LOGIC_VECTOR (31 downto 0));
end data_memory;

architecture Behavioral of data_memory is
type memory_file is array (0 to 258) of std_logic_vector (7 downto 0);
signal memory_data : memory_file:= (others => x"FF") ;
begin
process(clk) begin
    if(rising_edge(clk)) then
        if(wr_en ='1') then
            memory_data(to_integer(unsigned(addr))) <= wr_data(7 downto 0);
            memory_data(to_integer(unsigned(addr) +1)) <= wr_data(15 downto 8);
            memory_data(to_integer(unsigned(addr) +2)) <= wr_data(23 downto 16);
            memory_data(to_integer(unsigned(addr) +3)) <= wr_data(31 downto 24);
        end if;
    end if;
end process;
rd_data ( 7 downto 0) <= memory_data(to_integer(unsigned(addr)));
rd_data ( 15 downto 8) <= memory_data(to_integer(unsigned(addr)+1));
rd_data ( 23 downto 16) <= memory_data(to_integer(unsigned(addr)+2));
rd_data ( 31 downto 24) <= memory_data(to_integer(unsigned(addr)+3));

end Behavioral;